LIBRARY ieee ;
USE ieee.std_logic_1164.all ;

ENTITY guette_le_cpu IS
	PORT(
		


	);
END guette_le_cpu;



